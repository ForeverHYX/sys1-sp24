`ifdef VERILATE
    localparam FILE_PATH="initial.hex";
`else
    localparam FILE_PATH=;//your initial.hex
`endif