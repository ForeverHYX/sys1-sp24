`define DISPLAY 128'h01234567_89abcdef_00000032_30102930
//replace xxxxxx with your student ID