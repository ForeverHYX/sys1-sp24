module FSM(
    input rstn,
    input clk,
    input a,
    input b,
    output [1:0] state
);

    // fill your code

endmodule