module main( 
   input I0,
   input I1,
   input I2,
   input I3,
   output O 
);

   //your verilog code
   
endmodule
