module top(
  input SW0,
  input SW1,
  input SW2,
  input SW3,
  output LD0
);

  // add connection from FPGA IO to the main

endmodule