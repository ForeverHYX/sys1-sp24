/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : logisimTopLevelShell                                         **
 **                                                                          **
 *****************************************************************************/

module logisimTopLevelShell(  );

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire       s_I0;
   wire       s_I1;
   wire       s_I2;
   wire       s_I3;
   wire       s_O;
   wire [1:0] s_S;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** All signal adaptations are performed here                                  **
   *******************************************************************************/
   assign s_I0   = 1'b0;
   assign s_I1   = 1'b0;
   assign s_I2   = 1'b0;
   assign s_I3   = 1'b0;
   assign s_S[0] = 1'b0;
   assign s_S[1] = 1'b0;

   /*******************************************************************************
   ** The toplevel component is connected here                                   **
   *******************************************************************************/
   MUX4T1_1   CIRCUIT_0 (.I0(s_I0),
                         .I1(s_I1),
                         .I2(s_I2),
                         .I3(s_I3),
                         .O(s_O),
                         .S(s_S));
endmodule
